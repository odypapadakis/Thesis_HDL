`timescale 1ns / 1ns   // <time_unit> / <time_precision>


module Pseudo_Memory;






endmodule